module part1 (PIN_N2, PIN_G26);
  input PIN_N2, PIN_G26;

  //nios_system CPU (PIN_N2, DMAtS, DMB, DMD, DMR, DMWR, DMW, DMWD, IMAtS, IMR, JDMRD, JDMRR, PIN_G26, DMGJDM, DMQRJDM, DMRDVJDM, DMRJDM, IMGJDM, IMQRJDM, IMRDVJDM, JDMA, JDMBT, JDMB, JDMCS, JDMDA, JDMRDfSA, JDMRn, JDMRRfSA, JDMW, JDMWD, JDMEX)
  nios_system CPU0 (PIN_N2, PIN_G26);

endmodule
